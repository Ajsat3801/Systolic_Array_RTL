module instr_buffer #(

)(
    input clk,
    input [63:0] interface_input,
    output reg [63:0] instr_to_controller
)
endmodule